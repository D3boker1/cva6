/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
module bootrom_64 (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic [63:0]  addr_i,
   output logic [63:0]  rdata_o
);
    localparam int RomSize = 998;

    const logic [RomSize-1:0][63:0] mem = {
        64'h00000000_00000000,
        64'h0a0d2165_6e6f6420,
        64'h00000000_00206567,
        64'h616d6920_746f6f62,
        64'h20676e69_79706f63,
        64'h00000000_00000009,
        64'h3a656d61_6e090a0d,
        64'h00093a73_65747562,
        64'h69727474_61090a0d,
        64'h00000009_3a61626c,
        64'h20747361_6c090a0d,
        64'h0000093a_61626c20,
        64'h74737269_66090a0d,
        64'h00000000_00000000,
        64'h09202020_20203a64,
        64'h69756720_6e6f6974,
        64'h69747261_70090a0d,
        64'h00000000_00000000,
        64'h093a6469_75672065,
        64'h70797420_6e6f6974,
        64'h69747261_70090a0d,
        64'h00000000_20797274,
        64'h6e65206e_6f697469,
        64'h74726170_20747067,
        64'h00000009_20203a73,
        64'h65697274_6e65206e,
        64'h6f697469_74726170,
        64'h20657a69_73090a0d,
        64'h00000009_3a736569,
        64'h72746e65_206e6f69,
        64'h74697472_61702072,
        64'h65626d75_6e090a0d,
        64'h00000009_2020203a,
        64'h61626c20_73656972,
        64'h746e6520_6e6f6974,
        64'h69747261_70090a0d,
        64'h00093a61_646c2070,
        64'h756b6361_62090a0d,
        64'h00000000_00000000,
        64'h093a6162_6c20746e,
        64'h65727275_63090a0d,
        64'h00000009_3a646576,
        64'h72657365_72090a0d,
        64'h00093a72_65646165,
        64'h685f6372_63090a0d,
        64'h00000000_00000909,
        64'h3a657a69_73090a0d,
        64'h00000009_3a6e6f69,
        64'h73697665_72090a0d,
        64'h0000093a_65727574,
        64'h616e6769_73090a0d,
        64'h00000000_003a7265,
        64'h64616568_20656c62,
        64'h6174206e_6f697469,
        64'h74726170_20747067,
        64'h0000203a_65756c61,
        64'h76206e72_75746572,
        64'h2079706f_63206473,
        64'h00000000_0000000a,
        64'h0d216465_6c696166,
        64'h20647261_63204453,
        64'h00000000_0000000a,
        64'h0d216465_7a696c61,
        64'h6974696e_69206473,
        64'h00000000_0a0d676e,
        64'h69746978_65202e2e,
        64'h2e647320_657a696c,
        64'h61697469_6e692074,
        64'h6f6e2064_6c756f63,
        64'h00000000_0000002e,
        64'h00000000_0000000a,
        64'h0d6b636f_6c622044,
        64'h53206461_65722074,
        64'h6f6e2064_6c756f63,
        64'h0000000a_0d202e2e,
        64'h2e445320_676e697a,
        64'h696c6169_74696e69,
        64'h00000031_34646d63,
        64'h00000035_35646d63,
        64'h00000000_30646d63,
        64'h00000020_3a206573,
        64'h6e6f7073_65720920,
        64'h00000000_0020646e,
        64'h616d6d6f_63204453,
        64'h00000000_203f3f79,
        64'h74706d65_20746f6e,
        64'h206f6669_66207872,
        64'h00000000_00000a0d,
        64'h2164657a_696c6169,
        64'h74696e69_20495053,
        64'h00000000_00007830,
        64'h203a7375_74617473,
        64'h00000000_00000a0d,
        64'h49505320_74696e69,
        64'h00000a0d_21646c72,
        64'h6f57206f_6c6c6548,
        64'h00000000_00000032,
        64'h2d746c75_61666564,
        64'h2d697274_2c786e6c,
        64'h7800746c_75616665,
        64'h642d6972_742c786e,
        64'h6c78006c_6175642d,
        64'h73692c78_6e6c7800,
        64'h746e6573_6572702d,
        64'h74707572_7265746e,
        64'h692c786e_6c780068,
        64'h74646977_2d326f69,
        64'h70672c78_6e6c7800,
        64'h68746469_772d6f69,
        64'h70672c78_6e6c7800,
        64'h322d746c_75616665,
        64'h642d7475_6f642c78,
        64'h6e6c7800_746c7561,
        64'h6665642d_74756f64,
        64'h2c786e6c_7800322d,
        64'h73747570_6e692d6c,
        64'h6c612c78_6e6c7800,
        64'h73747570_6e692d6c,
        64'h6c612c78_6e6c7800,
        64'h72656c6c_6f72746e,
        64'h6f632d6f_69706700,
        64'h736c6c65_632d6f69,
        64'h70672300_73736572,
        64'h6464612d_63616d2d,
        64'h6c61636f_6c007077,
        64'h2d656c62_61736964,
        64'h00736567_6e61722d,
        64'h65676174_6c6f7600,
        64'h79636e65_75716572,
        64'h662d7861_6d2d6970,
        64'h73006f69_7461722d,
        64'h6b63732c_786e6c78,
        64'h00737469_622d7265,
        64'h66736e61_72742d6d,
        64'h756e2c78_6e6c7800,
        64'h73746962_2d73732d,
        64'h6d756e2c_786e6c78,
        64'h00747369_78652d6f,
        64'h6669662c_786e6c78,
        64'h00796c69_6d61662c,
        64'h786e6c78_00687464,
        64'h69772d6f_692d6765,
        64'h72007466_6968732d,
        64'h67657200_73747075,
        64'h72726574_6e690074,
        64'h6e657261_702d7470,
        64'h75727265_746e6900,
        64'h64656570_732d746e,
        64'h65727275_63007665,
        64'h646e2c76_63736972,
        64'h00797469_726f6972,
        64'h702d7861_6d2c7663,
        64'h73697200_73656d61,
        64'h6e2d6765_72006465,
        64'h646e6574_78652d73,
        64'h74707572_7265746e,
        64'h69007365_676e6172,
        64'h00646564_6e657073,
        64'h75732d65_74617473,
        64'h2d6e6961_74657200,
        64'h72656767_6972742d,
        64'h746c7561_6665642c,
        64'h78756e69_6c00736f,
        64'h69706700_656c646e,
        64'h61687000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h00736c6c_65632d74,
        64'h70757272_65746e69,
        64'h23007469_6c70732d,
        64'h626c7400_65707974,
        64'h2d756d6d_00617369,
        64'h2c766373_69720073,
        64'h75746174_73006765,
        64'h72006570_79745f65,
        64'h63697665_64007963,
        64'h6e657571_6572662d,
        64'h6b636f6c_63007963,
        64'h6e657571_6572662d,
        64'h65736162_656d6974,
        64'h00687461_702d7475,
        64'h6f647473_006c6564,
        64'h6f6d0065_6c626974,
        64'h61706d6f_6300736c,
        64'h6c65632d_657a6973,
        64'h2300736c_6c65632d,
        64'h73736572_64646123,
        64'h09000000_02000000,
        64'h02000000_02000000,
        64'h01000000_b5000000,
        64'h04000000_03000000,
        64'hffffffff_bf020000,
        64'h04000000_03000000,
        64'hffffffff_ae020000,
        64'h04000000_03000000,
        64'h01000000_a1020000,
        64'h04000000_03000000,
        64'h00000000_8a020000,
        64'h04000000_03000000,
        64'h08000000_79020000,
        64'h04000000_03000000,
        64'h08000000_69020000,
        64'h04000000_03000000,
        64'h00000000_55020000,
        64'h04000000_03000000,
        64'h00000000_43020000,
        64'h04000000_03000000,
        64'h00000000_31020000,
        64'h04000000_03000000,
        64'h00000000_21020000,
        64'h04000000_03000000,
        64'h00000100_00000000,
        64'h00000040_00000000,
        64'h67000000_10000000,
        64'h03000000_11020000,
        64'h00000000_03000000,
        64'h00000000_612e3030,
        64'h2e312d6f_6970672d,
        64'h7370782c_786e6c78,
        64'h1b000000_15000000,
        64'h03000000_02000000,
        64'h05020000_04000000,
        64'h03000000_00000030,
        64'h30303030_30303440,
        64'h6f697067_01000000,
        64'h02000000_00800000,
        64'h00000000_00000030,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h00007fe3_023e1800,
        64'hf3010000_06000000,
        64'h03000000_00000000,
        64'h03000000_52010000,
        64'h08000000_03000000,
        64'h04000000_41010000,
        64'h04000000_03000000,
        64'h006b726f_7774656e,
        64'h5b000000_08000000,
        64'h03000000_00687465,
        64'h2d637369_72776f6c,
        64'h1b000000_0c000000,
        64'h03000000_00000000,
        64'h30303030_30303033,
        64'h40687465_2d637369,
        64'h72776f6c_01000000,
        64'h02000000_02000000,
        64'he8010000_00000000,
        64'h03000000_e40c0000,
        64'he40c0000_d9010000,
        64'h08000000_03000000,
        64'h20bcbe00_c7010000,
        64'h04000000_03000000,
        64'h00000000_67000000,
        64'h04000000_03000000,
        64'h00000000_746f6c73,
        64'h2d697073_2d636d6d,
        64'h1b000000_0d000000,
        64'h03000000_00000030,
        64'h40636d6d_01000000,
        64'h04000000_b8010000,
        64'h04000000_03000000,
        64'h08000000_a1010000,
        64'h04000000_03000000,
        64'h01000000_90010000,
        64'h04000000_03000000,
        64'h01000000_80010000,
        64'h04000000_03000000,
        64'h00377865_746e696b,
        64'h74010000_08000000,
        64'h03000000_00100000,
        64'h00000000_00000020,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h02000000_02000000,
        64'h52010000_08000000,
        64'h03000000_04000000,
        64'h41010000_04000000,
        64'h03000000_00000000,
        64'h0f000000_04000000,
        64'h03000000_01000000,
        64'h00000000_04000000,
        64'h03000000_00612e30,
        64'h302e322d_6970732d,
        64'h7370782c_786e6c78,
        64'h00622e30_302e322d,
        64'h6970732d_7370782c,
        64'h786e6c78_1b000000,
        64'h28000000_03000000,
        64'h00000000_30303030,
        64'h30303032_40697073,
        64'h2d737078_01000000,
        64'h02000000_006c6f72,
        64'h746e6f63_0b010000,
        64'h08000000_03000000,
        64'h04000000_41010000,
        64'h04000000_03000000,
        64'h00100000_00000000,
        64'h00000018_00000000,
        64'h67000000_10000000,
        64'h03000000_07000000,
        64'h06000000_05000000,
        64'h04000000_52010000,
        64'h10000000_03000000,
        64'h00007265_6d69745f,
        64'h6270612c_706c7570,
        64'h1b000000_0f000000,
        64'h03000000_00003030,
        64'h30303030_38314072,
        64'h656d6974_01000000,
        64'h02000000_04000000,
        64'h67010000_04000000,
        64'h03000000_02000000,
        64'h5d010000_04000000,
        64'h03000000_01000000,
        64'h52010000_04000000,
        64'h03000000_04000000,
        64'h41010000_04000000,
        64'h03000000_00c20100,
        64'h33010000_04000000,
        64'h03000000_80f0fa02,
        64'h4b000000_04000000,
        64'h03000000_00100000,
        64'h00000000_00000010,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h00000000_61303535,
        64'h3631736e_1b000000,
        64'h09000000_03000000,
        64'h00000030_30303030,
        64'h30303140_74726175,
        64'h01000000_02000000,
        64'h04000000_b5000000,
        64'h04000000_03000000,
        64'h1e000000_28010000,
        64'h04000000_03000000,
        64'h07000000_15010000,
        64'h04000000_03000000,
        64'h00000004_00000000,
        64'h0000000c_00000000,
        64'h67000000_10000000,
        64'h03000000_09000000,
        64'h03000000_0b000000,
        64'h03000000_09000000,
        64'h02000000_0b000000,
        64'h02000000_f7000000,
        64'h20000000_03000000,
        64'ha0000000_00000000,
        64'h03000000_00306369,
        64'h6c702c76_63736972,
        64'h1b000000_0c000000,
        64'h03000000_01000000,
        64'h8f000000_04000000,
        64'h03000000_00000000,
        64'h00000000_04000000,
        64'h03000000_00000000,
        64'h30303030_30306340,
        64'h72656c6c_6f72746e,
        64'h6f632d74_70757272,
        64'h65746e69_01000000,
        64'h02000000_006c6f72,
        64'h746e6f63_0b010000,
        64'h08000000_03000000,
        64'h00000c00_00000000,
        64'h00000002_00000000,
        64'h67000000_10000000,
        64'h03000000_07000000,
        64'h03000000_03000000,
        64'h03000000_07000000,
        64'h02000000_03000000,
        64'h02000000_f7000000,
        64'h20000000_03000000,
        64'h00000000_30746e69,
        64'h6c632c76_63736972,
        64'h1b000000_0d000000,
        64'h03000000_00000030,
        64'h30303030_30324074,
        64'h6e696c63_01000000,
        64'hf0000000_00000000,
        64'h03000000_00007375,
        64'h622d656c_706d6973,
        64'h00636f73_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h1f000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00636f73_01000000,
        64'h02000000_02000000,
        64'hd9000000_00000000,
        64'h03000000_00000074,
        64'h61656274_72616568,
        64'hc3000000_0a000000,
        64'h03000000_00000000,
        64'h01000000_01000000,
        64'hbd000000_0c000000,
        64'h03000000_00000064,
        64'h656c2d74_61656274,
        64'h72616568_01000000,
        64'h00000073_64656c2d,
        64'h6f697067_1b000000,
        64'h0a000000_03000000,
        64'h00000000_7364656c,
        64'h01000000_02000000,
        64'h00000040_00000000,
        64'h00000080_00000000,
        64'h67000000_10000000,
        64'h03000000_00007972,
        64'h6f6d656d_5b000000,
        64'h07000000_03000000,
        64'h00303030_30303030,
        64'h38407972_6f6d656d,
        64'h01000000_02000000,
        64'h02000000_02000000,
        64'h03000000_b5000000,
        64'h04000000_03000000,
        64'h00006374_6e692d75,
        64'h70632c76_63736972,
        64'h1b000000_0f000000,
        64'h03000000_a0000000,
        64'h00000000_03000000,
        64'h01000000_8f000000,
        64'h04000000_03000000,
        64'h00000000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h01000000_85000000,
        64'h00000000_03000000,
        64'h00003933_76732c76,
        64'h63736972_7c000000,
        64'h0b000000_03000000,
        64'h00006364_66616d69,
        64'h34367672_72000000,
        64'h0b000000_03000000,
        64'h00000076_63736972,
        64'h00656e61_69726120,
        64'h2c687465_1b000000,
        64'h12000000_03000000,
        64'h00000000_79616b6f,
        64'h6b000000_05000000,
        64'h03000000_01000000,
        64'h67000000_04000000,
        64'h03000000_00757063,
        64'h5b000000_04000000,
        64'h03000000_005a6202,
        64'h4b000000_04000000,
        64'h03000000_00000031,
        64'h40757063_01000000,
        64'h02000000_02000000,
        64'h02000000_b5000000,
        64'h04000000_03000000,
        64'h00006374_6e692d75,
        64'h70632c76_63736972,
        64'h1b000000_0f000000,
        64'h03000000_a0000000,
        64'h00000000_03000000,
        64'h01000000_8f000000,
        64'h04000000_03000000,
        64'h00000000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h01000000_85000000,
        64'h00000000_03000000,
        64'h00003933_76732c76,
        64'h63736972_7c000000,
        64'h0b000000_03000000,
        64'h00006364_66616d69,
        64'h34367672_72000000,
        64'h0b000000_03000000,
        64'h00000076_63736972,
        64'h00656e61_69726120,
        64'h2c687465_1b000000,
        64'h12000000_03000000,
        64'h00000000_79616b6f,
        64'h6b000000_05000000,
        64'h03000000_00000000,
        64'h67000000_04000000,
        64'h03000000_00757063,
        64'h5b000000_04000000,
        64'h03000000_005a6202,
        64'h4b000000_04000000,
        64'h03000000_00000030,
        64'h40757063_01000000,
        64'h002d3101_38000000,
        64'h04000000_03000000,
        64'h00000000_0f000000,
        64'h04000000_03000000,
        64'h01000000_00000000,
        64'h04000000_03000000,
        64'h00000000_73757063,
        64'h01000000_02000000,
        64'h00000030_30323531,
        64'h313a3030_30303030,
        64'h30314074_7261752f,
        64'h636f732f_2c000000,
        64'h1a000000_03000000,
        64'h00006e65_736f6863,
        64'h01000000_00657261,
        64'h622d656e_61697261,
        64'h2c687465_26000000,
        64'h10000000_03000000,
        64'h00766564_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h14000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00000000_01000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h200a0000_d2020000,
        64'h00000000_10000000,
        64'h11000000_28000000,
        64'h580a0000_38000000,
        64'h2a0d0000_edfe0dd0,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h46454443_42413938,
        64'h37363534_33323130,
        64'h00000000_00000000,
        64'h00000000_00008067,
        64'h01010113_00000513,
        64'h00813083_c75ff0ef,
        64'h01f51513_000085b7,
        64'h00100513_bb4ff0ef,
        64'he6850513_00001517,
        64'hb78ff0ef_00113423,
        64'ha0050513_20058593,
        64'hff010113_02626537,
        64'h0001c5b7_cf9ff06f,
        64'hbe0ff0ef_18450513,
        64'h00001517_d95ff06f,
        64'hee050513_00001517,
        64'hcb8ff0ef_00090513,
        64'hc00ff0ef_fe450513,
        64'h00001517_c0cff0ef,
        64'hfd850513_00001517,
        64'hdc1ff06f_f0c50513,
        64'h00001517_ce4ff0ef,
        64'h00048513_c2cff0ef,
        64'h01050513_00001517,
        64'hc38ff0ef_00450513,
        64'h00001517_04050e63,
        64'h00050493_b5dff0ef,
        64'h40b6063b_0016061b,
        64'h000a0513_020aa583,
        64'h028ab603_c64ff0ef,
        64'h1f050513_00001517,
        64'hf36918e3_08048493,
        64'hc78ff0ef_0019091b,
        64'hf7050513_00001517,
        64'hff899ae3_dacff0ef,
        64'h00198993_0009c503,
        64'hc98ff0ef_21450513,
        64'h00001517_d64ff0ef,
        64'h0104b503_cacff0ef,
        64'h21850513_00001517,
        64'hd78ff0ef_0084b503,
        64'hcc0ff0ef_21c50513,
        64'h00001517_d8cff0ef,
        64'h06048c13_01848993,
        64'h0004b503_cdcff0ef,
        64'h22850513_00001517,
        64'hff349ae3_e0cff0ef,
        64'h00198993_0009c503,
        64'hff048993_cfcff0ef,
        64'h22850513_00001517,
        64'hff7998e3_e2cff0ef,
        64'h00198993_0007c503,
        64'h013c07b3_00000993,
        64'hd20ff0ef_fe048c13,
        64'h23050513_00001517,
        64'he50ff0ef_0ff97513,
        64'hd38ff0ef_22c50513,
        64'h00001517_00400b13,
        64'h01000b93_12051c63,
        64'h02010493_00050913,
        64'h00010a93_c6dff0ef,
        64'h00010513_00100613,
        64'he0010113_04892583,
        64'hd70ff0ef_06450513,
        64'h00001517_ddcff0ef,
        64'h05412503_d84ff0ef,
        64'h25850513_00001517,
        64'hdf0ff0ef_05012503,
        64'hd98ff0ef_24c50513,
        64'h00001517_e64ff0ef,
        64'h04813503_dacff0ef,
        64'h24050513_00001517,
        64'he78ff0ef_02013503,
        64'hdc0ff0ef_24450513,
        64'h00001517_e8cff0ef,
        64'h01813503_dd4ff0ef,
        64'h24050513_00001517,
        64'he40ff0ef_01412503,
        64'hde8ff0ef_24450513,
        64'h00001517_e54ff0ef,
        64'h01012503_dfcff0ef,
        64'h24850513_00001517,
        64'he68ff0ef_00c12503,
        64'he10ff0ef_24c50513,
        64'h00001517_e7cff0ef,
        64'h00812503_e24ff0ef,
        64'h25050513_00001517,
        64'hef0ff0ef_00013503,
        64'he38ff0ef_25450513,
        64'h00001517_e44ff0ef,
        64'h24050513_00001517,
        64'hf6dff06f_ffe00493,
        64'he58ff0ef_14c50513,
        64'h00001517_f24ff0ef,
        64'h00048513_e6cff0ef,
        64'h25050513_00001517,
        64'he78ff0ef_24450513,
        64'h00001517_02050c63,
        64'h00050493_00010913,
        64'hda1ff0ef_00010513,
        64'h00100593_00100613,
        64'he0010113_ea4ff0ef,
        64'h25850513_00001517,
        64'h00008067_05010113,
        64'h00013c03_00813b83,
        64'h01013b03_01813a83,
        64'h02013a03_02813983,
        64'h03013903_03813483,
        64'h04013403_00048513,
        64'h04813083_fb040113,
        64'hfff00493_eecff0ef,
        64'h27850513_00001517,
        64'h04050663_d25ff0ef,
        64'h00050a13_05010413,
        64'h01813023_01713423,
        64'h01613823_01513c23,
        64'h03313423_03213823,
        64'h02913c23_04113423,
        64'h03413023_04813023,
        64'hfb010113_f85ff06f,
        64'hffe00413_00008067,
        64'h0d010113_08813b83,
        64'h09013b03_09813a83,
        64'h0a013a03_0a813983,
        64'h0b013903_0b813483,
        64'h0c013403_00040513,
        64'h0c813083_fff00413,
        64'hf70ff0ef_2d450513,
        64'h00001517_b09ff0ef,
        64'hb0dff0ef_b11ff0ef,
        64'hb15ff0ef_b19ff0ef,
        64'hb1dff0ef_b21ff0ef,
        64'hb25ff0ef_0340006f,
        64'hb2dff0ef_b39ff0ef,
        64'h00c00513_00000593,
        64'h00100613_00000413,
        64'hf72046e3_fff90913,
        64'hfc0ff0ef_34450513,
        64'h00001517_00079863,
        64'h034967b3_08941e63,
        64'h0004849b_03045413,
        64'h03041413_00a46433,
        64'hb75ff0ef_03045413,
        64'h03041413_0085141b,
        64'h00040a93_b89ff0ef,
        64'hfd6414e3_04040413,
        64'hff7a94e3_00050493,
        64'hecdff0ef_001a8a93,
        64'h00048513_0007c583,
        64'h015407b3_04000b93,
        64'h00000a93_b01ff0ef,
        64'h00010513_04000593,
        64'h00040613_200a8b13,
        64'h00000493_000a8413,
        64'hff351ee3_bd9ff0ef,
        64'h3e800a13_0fe00993,
        64'h0c051063_bf1ff0ef,
        64'h01200513_00040593,
        64'h0ff67613_00166613,
        64'h0015161b_f05ff0ef,
        64'h0ff47593_f0dff0ef,
        64'h0ff5f593_0084559b,
        64'hf19ff0ef_0ff5f593,
        64'h0104559b_f25ff0ef,
        64'h00000513_0184559b,
        64'hfee79ae3_00178793,
        64'h00c68023_00f106b3,
        64'h08000713_fff00613,
        64'h00000793_02095913,
        64'h00058413_00050a93,
        64'h09713423_09613823,
        64'h0b413023_0b313423,
        64'h0a913c23_0c113423,
        64'h09513c23_0c813023,
        64'h02061913_0b213823,
        64'hf3010113_00008067,
        64'h03055513_03051513,
        64'h00f54533_00e7f7b3,
        64'hfe078793_0057171b,
        64'h000027b7_0107571b,
        64'h0105171b_00f54533,
        64'h00c5179b_00b54533,
        64'h00f57513_0045d51b,
        64'h00b7c5b3_0307d793,
        64'h03079793_00a7e7b3,
        64'h0085551b_0085179b,
        64'h00008067_07f57513,
        64'h00f54533_0ff7f793,
        64'h0045179b_00b54533,
        64'h0ff57513_00f54533,
        64'h0045d51b_0075d79b,
        64'h00b575b3_00008067,
        64'h01010113_00078513,
        64'h00013403_00813083,
        64'hffd00793_00051463,
        64'h00000793_f5dff0ef,
        64'h00050a63_ffe00793,
        64'he99ff0ef_02050063,
        64'hfff00793_e2dff0ef,
        64'hfe041ce3_d41ff0ef,
        64'hfff4041b_00a00413,
        64'h9c1ff0ef_50c50513,
        64'h00001517_b25ff0ef,
        64'h00813023_00113423,
        64'hff010113_00008067,
        64'h02010113_00153513,
        64'h00813483_01013403,
        64'h0004051b_01813083,
        64'hfc940ae3_d89ff0ef,
        64'he25ff0ef_54450513,
        64'h00001517_00050593,
        64'h00050413_da9ff0ef,
        64'h02900513_400005b7,
        64'h07700613_f9dff0ef,
        64'h00100493_00813823,
        64'h00113c23_00913423,
        64'hfe010113_00008067,
        64'h01010113_00153513,
        64'hfff50513_00013403,
        64'h0004051b_00813083,
        64'he7dff0ef_59850513,
        64'h00040593_00001517,
        64'hdf5ff0ef_00050413,
        64'he05ff0ef_00813023,
        64'h00113423_03700513,
        64'h00000593_06500613,
        64'hff010113_00008067,
        64'h02010113_00013903,
        64'h00813483_01013403,
        64'h01813083_00143513,
        64'hf5640413_0004041b,
        64'h01249863_00f4f493,
        64'h00f91c63_00000513,
        64'h00100793_e51ff0ef,
        64'he55ff0ef_00050413,
        64'he5dff0ef_00050493,
        64'he65ff0ef_e69ff0ef,
        64'he6dff0ef_00050913,
        64'he7dff0ef_01213023,
        64'h00913423_00813823,
        64'h00113c23_00800513,
        64'h1aa00593_08700613,
        64'hfe010113_fe5ff06f,
        64'h00000513_00008067,
        64'h02010113_00013903,
        64'h00813483_01013403,
        64'h01813083_00100513,
        64'hf55ff0ef_00100593,
        64'h66850513_00001517,
        64'hff2490e3_02040a63,
        64'hed5ff0ef_00050493,
        64'hfff4041b_ee9ff0ef,
        64'h00000513_00000593,
        64'h09500613_00100913,
        64'h71040413_00913423,
        64'h00113c23_01213023,
        64'h00002437_00813823,
        64'hfe010113_b85ff06f,
        64'h02010113_67c50513,
        64'h00001517_00813483,
        64'h01813083_01013403,
        64'hcc1ff0ef_00040513,
        64'hba9ff0ef_6cc50513,
        64'h00001517_bb5ff0ef,
        64'h00048513_bbdff0ef,
        64'h00058413_00813823,
        64'h00113c23_6dc50513,
        64'h00001517_00050493,
        64'h00913423_fe010113,
        64'h00008067_02010113,
        64'h00013903_00813483,
        64'h01013403_01813083,
        64'hfe0416e3_fff40413,
        64'h0007d663_4187d79b,
        64'h0185179b_f99ff0ef,
        64'h06400413_e35ff0ef,
        64'h00048513_e3dff0ef,
        64'h0ff47513_e45ff0ef,
        64'h0ff57513_0084551b,
        64'he51ff0ef_0ff57513,
        64'h0104551b_e5dff0ef,
        64'h0184551b_e65ff0ef,
        64'h04096513_fd9ff0ef,
        64'h00050913_01213023,
        64'h00060493_00058413,
        64'h00913423_00813823,
        64'h00113c23_fe010113,
        64'he91ff06f_0ff00513,
        64'h00008067_fff00513,
        64'hfadff06f_00d70023,
        64'h00178793_00f60733,
        64'h06c82683_fc0712e3,
        64'h00177713_06452703,
        64'hf91ff06f_06e6a423,
        64'h00178793_00074703,
        64'h00f50733_00008067,
        64'h00000513_06e7a023,
        64'h00600713_06e7a823,
        64'hfff00713_200007b7,
        64'h02b6ea63_0007869b,
        64'h20000837_20000537,
        64'hfe079ce3_0017f793,
        64'h06472783_20000737,
        64'h06e7a023_200007b7,
        64'h10600713_fe079ce3,
        64'hfff7879b_00000013,
        64'h03200793_04b76e63,
        64'h0007871b_00000793,
        64'h200006b7_06e7a823,
        64'hffe00713_200007b7,
        64'h0ab7e663_10000793,
        64'h00008067_02010113,
        64'h00813483_06e7a023,
        64'h00600713_06e7a823,
        64'h01013403_0ff47513,
        64'hfff00713_200007b7,
        64'h01813083_d5dff0ef,
        64'h85050513_00002517,
        64'he29ff0ef_02055513,
        64'h02051513_0004a503,
        64'hd79ff0ef_87450513,
        64'h00002517_02079663,
        64'h0017f793_0004041b,
        64'h0647a783_06c7a403,
        64'hfe071ae3_00177713,
        64'h06478493_0647a703,
        64'h06e7a023_10600713,
        64'h200007b7_fe079ce3,
        64'hfff7879b_00000013,
        64'h06400793_06a7a423,
        64'h06e7a823_ffe00713,
        64'h00913423_00813823,
        64'h00113c23_200007b7,
        64'hfe010113_de5ff06f,
        64'h02010113_8cc50513,
        64'h00002517_00813483,
        64'h01813083_01013403,
        64'h06f42023_00600793,
        64'he09ff0ef_8fc50513,
        64'h00002517_ed5ff0ef,
        64'h02055513_02049513,
        64'h0004849b_e25ff0ef,
        64'h8f850513_00002517,
        64'h06442483_06f42023,
        64'h16600793_e3dff0ef,
        64'h93050513_00002517,
        64'hf09ff0ef_02055513,
        64'h02049513_0004849b,
        64'he59ff0ef_92c50513,
        64'h00002517_06442483,
        64'h06f42023_10400793,
        64'h20000437_fe079ce3,
        64'hfff7879b_00000013,
        64'h00a00793_04e7a023,
        64'h00a00713_200007b7,
        64'he91ff0ef_00913423,
        64'h00813823_00113c23,
        64'h96450513_fe010113,
        64'h00002517_00008067,
        64'h00052503_00008067,
        64'h00b52023_e5dff06f,
        64'h02010113_01813083,
        64'h00914503_e6dff0ef,
        64'h00814503_f09ff0ef,
        64'h00113c23_00810593,
        64'hfe010113_00008067,
        64'h03010113_01013903,
        64'h01813483_02013403,
        64'h02813083_fd241ee3,
        64'hea1ff0ef_00914503,
        64'hea9ff0ef_ff84041b,
        64'h00814503_f49ff0ef,
        64'h0ff57513_00810593,
        64'h0084d533_ff800913,
        64'h03800413_00050493,
        64'h02113423_01213823,
        64'h00913c23_02813023,
        64'hfd010113_00008067,
        64'h03010113_01013903,
        64'h01813483_02013403,
        64'h02813083_fd241ee3,
        64'hf01ff0ef_00914503,
        64'hf09ff0ef_ff84041b,
        64'h00814503_fa9ff0ef,
        64'h0ff57513_00810593,
        64'h0084d53b_ff800913,
        64'h01800413_00050493,
        64'h02113423_01213823,
        64'h00913c23_02813023,
        64'hfd010113_00008067,
        64'h00f58023_0007c783,
        64'h00e580a3_00a787b3,
        64'h00455513_00074703,
        64'h00e78733_00f57713,
        64'hc4878793_00001797,
        64'hfe1ff06f_00140413,
        64'hf79ff0ef_00008067,
        64'h01010113_00013403,
        64'h00813083_00051a63,
        64'h00044503_00050413,
        64'h00113423_00813023,
        64'hff010113_00008067,
        64'h00e78823_02000713,
        64'h00e78423_fc700713,
        64'h00e78623_00300713,
        64'h00a78223_0ff57513,
        64'h00e78023_0085551b,
        64'h0ff57713_00e78623,
        64'hf8000713_00078223,
        64'h100007b7_02b5553b,
        64'h0045959b_00008067,
        64'h00a70023_fe078ce3,
        64'h0207f793_01474783,
        64'h10000737_00008067,
        64'h02057513_0147c503,
        64'h100007b7_00008067,
        64'h00054503_00008067,
        64'h00b50023_00008067,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00048067_01f49493,
        64'h0010049b_ea458593,
        64'h00001597_f1402573,
        64'h0924a4af_00190913,
        64'h04048493_01a49493,
        64'h0210049b_ff2496e3,
        64'hf14024f3_0004a903,
        64'h04048493_01a49493,
        64'h0210049b_585000ef,
        64'h01a11113_0210011b,
        64'h01249863_f1402973,
        64'h00000493_0924a4af,
        64'h00000913_04048493,
        64'h01a49493_0210049b
    };

    logic [$clog2(RomSize)-1:0] addr_q;

    always_ff @(posedge clk_i) begin
        if (req_i) begin
            addr_q <= addr_i[$clog2(RomSize)-1+3:3];
        end
    end

    // this prevents spurious Xes from propagating into
    // the speculative fetch stage of the core
    assign rdata_o = (addr_q < RomSize) ? mem[addr_q] : '0;
endmodule
