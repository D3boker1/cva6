/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
module bootrom_64 (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic [63:0]  addr_i,
   output logic [63:0]  rdata_o
);
    localparam int RomSize = 1030;

    const logic [RomSize-1:0][63:0] mem = {
        64'h00000000_00000000,
        64'h0a0d2165_6e6f6420,
        64'h00000000_00206567,
        64'h616d6920_746f6f62,
        64'h20676e69_79706f63,
        64'h00000000_00000009,
        64'h3a656d61_6e090a0d,
        64'h00093a73_65747562,
        64'h69727474_61090a0d,
        64'h00000009_3a61626c,
        64'h20747361_6c090a0d,
        64'h0000093a_61626c20,
        64'h74737269_66090a0d,
        64'h00000000_00000000,
        64'h09202020_20203a64,
        64'h69756720_6e6f6974,
        64'h69747261_70090a0d,
        64'h00000000_00000000,
        64'h093a6469_75672065,
        64'h70797420_6e6f6974,
        64'h69747261_70090a0d,
        64'h00000000_20797274,
        64'h6e65206e_6f697469,
        64'h74726170_20747067,
        64'h00000009_20203a73,
        64'h65697274_6e65206e,
        64'h6f697469_74726170,
        64'h20657a69_73090a0d,
        64'h00000009_3a736569,
        64'h72746e65_206e6f69,
        64'h74697472_61702072,
        64'h65626d75_6e090a0d,
        64'h00000009_2020203a,
        64'h61626c20_73656972,
        64'h746e6520_6e6f6974,
        64'h69747261_70090a0d,
        64'h00093a61_646c2070,
        64'h756b6361_62090a0d,
        64'h00000000_00000000,
        64'h093a6162_6c20746e,
        64'h65727275_63090a0d,
        64'h00000009_3a646576,
        64'h72657365_72090a0d,
        64'h00093a72_65646165,
        64'h685f6372_63090a0d,
        64'h00000000_00000909,
        64'h3a657a69_73090a0d,
        64'h00000009_3a6e6f69,
        64'h73697665_72090a0d,
        64'h0000093a_65727574,
        64'h616e6769_73090a0d,
        64'h00000000_003a7265,
        64'h64616568_20656c62,
        64'h6174206e_6f697469,
        64'h74726170_20747067,
        64'h0000203a_65756c61,
        64'h76206e72_75746572,
        64'h2079706f_63206473,
        64'h00000000_0000000a,
        64'h0d216465_6c696166,
        64'h20647261_63204453,
        64'h00000000_0000000a,
        64'h0d216465_7a696c61,
        64'h6974696e_69206473,
        64'h00000000_0a0d676e,
        64'h69746978_65202e2e,
        64'h2e647320_657a696c,
        64'h61697469_6e692074,
        64'h6f6e2064_6c756f63,
        64'h00000000_0000002e,
        64'h00000000_0000000a,
        64'h0d6b636f_6c622044,
        64'h53206461_65722074,
        64'h6f6e2064_6c756f63,
        64'h0000000a_0d202e2e,
        64'h2e445320_676e697a,
        64'h696c6169_74696e69,
        64'h00000031_34646d63,
        64'h00000035_35646d63,
        64'h00000000_30646d63,
        64'h00000020_3a206573,
        64'h6e6f7073_65720920,
        64'h00000000_0020646e,
        64'h616d6d6f_63204453,
        64'h00000000_203f3f79,
        64'h74706d65_20746f6e,
        64'h206f6669_66207872,
        64'h00000000_00000a0d,
        64'h2164657a_696c6169,
        64'h74696e69_20495053,
        64'h00000000_00007830,
        64'h203a7375_74617473,
        64'h00000000_00000a0d,
        64'h49505320_74696e69,
        64'h00000a0d_21646c72,
        64'h6f57206f_6c6c6548,
        64'h00000000_00000032,
        64'h2d746c75_61666564,
        64'h2d697274_2c786e6c,
        64'h7800746c_75616665,
        64'h642d6972_742c786e,
        64'h6c78006c_6175642d,
        64'h73692c78_6e6c7800,
        64'h746e6573_6572702d,
        64'h74707572_7265746e,
        64'h692c786e_6c780068,
        64'h74646977_2d326f69,
        64'h70672c78_6e6c7800,
        64'h68746469_772d6f69,
        64'h70672c78_6e6c7800,
        64'h322d746c_75616665,
        64'h642d7475_6f642c78,
        64'h6e6c7800_746c7561,
        64'h6665642d_74756f64,
        64'h2c786e6c_7800322d,
        64'h73747570_6e692d6c,
        64'h6c612c78_6e6c7800,
        64'h73747570_6e692d6c,
        64'h6c612c78_6e6c7800,
        64'h72656c6c_6f72746e,
        64'h6f632d6f_69706700,
        64'h736c6c65_632d6f69,
        64'h70672300_73736572,
        64'h6464612d_63616d2d,
        64'h6c61636f_6c007077,
        64'h2d656c62_61736964,
        64'h00736567_6e61722d,
        64'h65676174_6c6f7600,
        64'h79636e65_75716572,
        64'h662d7861_6d2d6970,
        64'h73006f69_7461722d,
        64'h6b63732c_786e6c78,
        64'h00737469_622d7265,
        64'h66736e61_72742d6d,
        64'h756e2c78_6e6c7800,
        64'h73746962_2d73732d,
        64'h6d756e2c_786e6c78,
        64'h00747369_78652d6f,
        64'h6669662c_786e6c78,
        64'h00796c69_6d61662c,
        64'h786e6c78_00687464,
        64'h69772d6f_692d6765,
        64'h72007466_6968732d,
        64'h67657200_73747075,
        64'h72726574_6e690074,
        64'h6e657261_702d7470,
        64'h75727265_746e6900,
        64'h64656570_732d746e,
        64'h65727275_63007665,
        64'h646e2c76_63736972,
        64'h00797469_726f6972,
        64'h702d7861_6d2c7663,
        64'h73697200_73656d61,
        64'h6e2d6765_72006465,
        64'h646e6574_78652d73,
        64'h74707572_7265746e,
        64'h69007365_676e6172,
        64'h00646564_6e657073,
        64'h75732d65_74617473,
        64'h2d6e6961_74657200,
        64'h72656767_6972742d,
        64'h746c7561_6665642c,
        64'h78756e69_6c00736f,
        64'h69706700_656c646e,
        64'h61687000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h00736c6c_65632d74,
        64'h70757272_65746e69,
        64'h23007469_6c70732d,
        64'h626c7400_65707974,
        64'h2d756d6d_00617369,
        64'h2c766373_69720073,
        64'h75746174_73006765,
        64'h72006570_79745f65,
        64'h63697665_64007963,
        64'h6e657571_6572662d,
        64'h6b636f6c_63007963,
        64'h6e657571_6572662d,
        64'h65736162_656d6974,
        64'h00687461_702d7475,
        64'h6f647473_006c6564,
        64'h6f6d0065_6c626974,
        64'h61706d6f_6300736c,
        64'h6c65632d_657a6973,
        64'h2300736c_6c65632d,
        64'h73736572_64646123,
        64'h09000000_02000000,
        64'h02000000_02000000,
        64'h01000000_b5000000,
        64'h04000000_03000000,
        64'hffffffff_bf020000,
        64'h04000000_03000000,
        64'hffffffff_ae020000,
        64'h04000000_03000000,
        64'h01000000_a1020000,
        64'h04000000_03000000,
        64'h00000000_8a020000,
        64'h04000000_03000000,
        64'h08000000_79020000,
        64'h04000000_03000000,
        64'h08000000_69020000,
        64'h04000000_03000000,
        64'h00000000_55020000,
        64'h04000000_03000000,
        64'h00000000_43020000,
        64'h04000000_03000000,
        64'h00000000_31020000,
        64'h04000000_03000000,
        64'h00000000_21020000,
        64'h04000000_03000000,
        64'h00000100_00000000,
        64'h00000040_00000000,
        64'h67000000_10000000,
        64'h03000000_11020000,
        64'h00000000_03000000,
        64'h00000000_612e3030,
        64'h2e312d6f_6970672d,
        64'h7370782c_786e6c78,
        64'h1b000000_15000000,
        64'h03000000_02000000,
        64'h05020000_04000000,
        64'h03000000_00000030,
        64'h30303030_30303440,
        64'h6f697067_01000000,
        64'h02000000_00800000,
        64'h00000000_00000030,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h00007fe3_023e1800,
        64'hf3010000_06000000,
        64'h03000000_00000000,
        64'h03000000_52010000,
        64'h08000000_03000000,
        64'h04000000_41010000,
        64'h04000000_03000000,
        64'h006b726f_7774656e,
        64'h5b000000_08000000,
        64'h03000000_00687465,
        64'h2d637369_72776f6c,
        64'h1b000000_0c000000,
        64'h03000000_00000000,
        64'h30303030_30303033,
        64'h40687465_2d637369,
        64'h72776f6c_01000000,
        64'h02000000_02000000,
        64'he8010000_00000000,
        64'h03000000_e40c0000,
        64'he40c0000_d9010000,
        64'h08000000_03000000,
        64'h20bcbe00_c7010000,
        64'h04000000_03000000,
        64'h00000000_67000000,
        64'h04000000_03000000,
        64'h00000000_746f6c73,
        64'h2d697073_2d636d6d,
        64'h1b000000_0d000000,
        64'h03000000_00000030,
        64'h40636d6d_01000000,
        64'h04000000_b8010000,
        64'h04000000_03000000,
        64'h08000000_a1010000,
        64'h04000000_03000000,
        64'h01000000_90010000,
        64'h04000000_03000000,
        64'h01000000_80010000,
        64'h04000000_03000000,
        64'h00377865_746e696b,
        64'h74010000_08000000,
        64'h03000000_00100000,
        64'h00000000_00000020,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h02000000_02000000,
        64'h52010000_08000000,
        64'h03000000_04000000,
        64'h41010000_04000000,
        64'h03000000_00000000,
        64'h0f000000_04000000,
        64'h03000000_01000000,
        64'h00000000_04000000,
        64'h03000000_00612e30,
        64'h302e322d_6970732d,
        64'h7370782c_786e6c78,
        64'h00622e30_302e322d,
        64'h6970732d_7370782c,
        64'h786e6c78_1b000000,
        64'h28000000_03000000,
        64'h00000000_30303030,
        64'h30303032_40697073,
        64'h2d737078_01000000,
        64'h02000000_006c6f72,
        64'h746e6f63_0b010000,
        64'h08000000_03000000,
        64'h04000000_41010000,
        64'h04000000_03000000,
        64'h00100000_00000000,
        64'h00000018_00000000,
        64'h67000000_10000000,
        64'h03000000_07000000,
        64'h06000000_05000000,
        64'h04000000_52010000,
        64'h10000000_03000000,
        64'h00007265_6d69745f,
        64'h6270612c_706c7570,
        64'h1b000000_0f000000,
        64'h03000000_00003030,
        64'h30303030_38314072,
        64'h656d6974_01000000,
        64'h02000000_04000000,
        64'h67010000_04000000,
        64'h03000000_02000000,
        64'h5d010000_04000000,
        64'h03000000_01000000,
        64'h52010000_04000000,
        64'h03000000_04000000,
        64'h41010000_04000000,
        64'h03000000_00c20100,
        64'h33010000_04000000,
        64'h03000000_80f0fa02,
        64'h4b000000_04000000,
        64'h03000000_00100000,
        64'h00000000_00000010,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h00000000_61303535,
        64'h3631736e_1b000000,
        64'h09000000_03000000,
        64'h00000030_30303030,
        64'h30303140_74726175,
        64'h01000000_02000000,
        64'h04000000_b5000000,
        64'h04000000_03000000,
        64'h1e000000_28010000,
        64'h04000000_03000000,
        64'h07000000_15010000,
        64'h04000000_03000000,
        64'h00000004_00000000,
        64'h0000000c_00000000,
        64'h67000000_10000000,
        64'h03000000_09000000,
        64'h03000000_0b000000,
        64'h03000000_09000000,
        64'h02000000_0b000000,
        64'h02000000_f7000000,
        64'h20000000_03000000,
        64'ha0000000_00000000,
        64'h03000000_00306369,
        64'h6c702c76_63736972,
        64'h1b000000_0c000000,
        64'h03000000_01000000,
        64'h8f000000_04000000,
        64'h03000000_00000000,
        64'h00000000_04000000,
        64'h03000000_00000000,
        64'h30303030_30306340,
        64'h72656c6c_6f72746e,
        64'h6f632d74_70757272,
        64'h65746e69_01000000,
        64'h02000000_006c6f72,
        64'h746e6f63_0b010000,
        64'h08000000_03000000,
        64'h00000c00_00000000,
        64'h00000002_00000000,
        64'h67000000_10000000,
        64'h03000000_07000000,
        64'h03000000_03000000,
        64'h03000000_07000000,
        64'h02000000_03000000,
        64'h02000000_f7000000,
        64'h20000000_03000000,
        64'h00000000_30746e69,
        64'h6c632c76_63736972,
        64'h1b000000_0d000000,
        64'h03000000_00000030,
        64'h30303030_30324074,
        64'h6e696c63_01000000,
        64'hf0000000_00000000,
        64'h03000000_00007375,
        64'h622d656c_706d6973,
        64'h00636f73_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h1f000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00636f73_01000000,
        64'h02000000_02000000,
        64'hd9000000_00000000,
        64'h03000000_00000074,
        64'h61656274_72616568,
        64'hc3000000_0a000000,
        64'h03000000_00000000,
        64'h01000000_01000000,
        64'hbd000000_0c000000,
        64'h03000000_00000064,
        64'h656c2d74_61656274,
        64'h72616568_01000000,
        64'h00000073_64656c2d,
        64'h6f697067_1b000000,
        64'h0a000000_03000000,
        64'h00000000_7364656c,
        64'h01000000_02000000,
        64'h00000040_00000000,
        64'h00000080_00000000,
        64'h67000000_10000000,
        64'h03000000_00007972,
        64'h6f6d656d_5b000000,
        64'h07000000_03000000,
        64'h00303030_30303030,
        64'h38407972_6f6d656d,
        64'h01000000_02000000,
        64'h02000000_02000000,
        64'h03000000_b5000000,
        64'h04000000_03000000,
        64'h00006374_6e692d75,
        64'h70632c76_63736972,
        64'h1b000000_0f000000,
        64'h03000000_a0000000,
        64'h00000000_03000000,
        64'h01000000_8f000000,
        64'h04000000_03000000,
        64'h00000000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h01000000_85000000,
        64'h00000000_03000000,
        64'h00003933_76732c76,
        64'h63736972_7c000000,
        64'h0b000000_03000000,
        64'h00006364_66616d69,
        64'h34367672_72000000,
        64'h0b000000_03000000,
        64'h00000076_63736972,
        64'h00656e61_69726120,
        64'h2c687465_1b000000,
        64'h12000000_03000000,
        64'h00000000_79616b6f,
        64'h6b000000_05000000,
        64'h03000000_01000000,
        64'h67000000_04000000,
        64'h03000000_00757063,
        64'h5b000000_04000000,
        64'h03000000_80f0fa02,
        64'h4b000000_04000000,
        64'h03000000_00000031,
        64'h40757063_01000000,
        64'h02000000_02000000,
        64'h02000000_b5000000,
        64'h04000000_03000000,
        64'h00006374_6e692d75,
        64'h70632c76_63736972,
        64'h1b000000_0f000000,
        64'h03000000_a0000000,
        64'h00000000_03000000,
        64'h01000000_8f000000,
        64'h04000000_03000000,
        64'h00000000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h01000000_85000000,
        64'h00000000_03000000,
        64'h00003933_76732c76,
        64'h63736972_7c000000,
        64'h0b000000_03000000,
        64'h00006364_66616d69,
        64'h34367672_72000000,
        64'h0b000000_03000000,
        64'h00000076_63736972,
        64'h00656e61_69726120,
        64'h2c687465_1b000000,
        64'h12000000_03000000,
        64'h00000000_79616b6f,
        64'h6b000000_05000000,
        64'h03000000_00000000,
        64'h67000000_04000000,
        64'h03000000_00757063,
        64'h5b000000_04000000,
        64'h03000000_80f0fa02,
        64'h4b000000_04000000,
        64'h03000000_00000030,
        64'h40757063_01000000,
        64'h40787d01_38000000,
        64'h04000000_03000000,
        64'h00000000_0f000000,
        64'h04000000_03000000,
        64'h01000000_00000000,
        64'h04000000_03000000,
        64'h00000000_73757063,
        64'h01000000_02000000,
        64'h00000030_30323531,
        64'h313a3030_30303030,
        64'h30314074_7261752f,
        64'h636f732f_2c000000,
        64'h1a000000_03000000,
        64'h00006e65_736f6863,
        64'h01000000_00657261,
        64'h622d656e_61697261,
        64'h2c687465_26000000,
        64'h10000000_03000000,
        64'h00766564_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h14000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00000000_01000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h200a0000_d2020000,
        64'h00000000_10000000,
        64'h11000000_28000000,
        64'h580a0000_38000000,
        64'h2a0d0000_edfe0dd0,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h46454443_42413938,
        64'h37363534_33323130,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00008067,
        64'h01010113_00000513,
        64'h00813083_c69ff0ef,
        64'h01f51513_000085b7,
        64'h00100513_ba0ff0ef,
        64'hf5050513_00001517,
        64'hb64ff0ef_00113423,
        64'h08050513_20058593,
        64'hff010113_02faf537,
        64'h0001c5b7_cf1ff06f,
        64'hbccff0ef_26c50513,
        64'h00001517_d91ff06f,
        64'hfc850513_00001517,
        64'hca4ff0ef_00048513,
        64'hbecff0ef_0cc50513,
        64'h00001517_bf8ff0ef,
        64'h0c050513_00001517,
        64'hdbdff06f_ff450513,
        64'h00001517_cd0ff0ef,
        64'h00048513_c18ff0ef,
        64'h0f850513_00001517,
        64'hc24ff0ef_0ec50513,
        64'h00001517_04050e63,
        64'h00050493_b4dff0ef,
        64'h40b6063b_0016061b,
        64'h000b0513_020aa583,
        64'h028ab603_c50ff0ef,
        64'h2d850513_00001517,
        64'hf37498e3_08090913,
        64'h080a0993_c68ff0ef,
        64'h0014849b_05c50513,
        64'h00001517_ff3a1ae3,
        64'hd9cff0ef_001a0a13,
        64'h000a4503_c88ff0ef,
        64'h30050513_00001517,
        64'hd54ff0ef_01093503,
        64'hc9cff0ef_30450513,
        64'h00001517_d68ff0ef,
        64'h00893503_cb0ff0ef,
        64'h30850513_00001517,
        64'hd7cff0ef_fb898a13,
        64'h00093503_cc8ff0ef,
        64'h31050513_00001517,
        64'hff2a1ae3_df8ff0ef,
        64'h001a0a13_000a4503,
        64'hf9098a13_ce8ff0ef,
        64'h31050513_00001517,
        64'hff8a18e3_e18ff0ef,
        64'h001a0a13_0007c503,
        64'h014c87b3_00000a13,
        64'hd0cff0ef_f8098c93,
        64'h31850513_00001517,
        64'he3cff0ef_0ff4f513,
        64'hd24ff0ef_31450513,
        64'h00001517_00400b93,
        64'h01000c13_12051c63,
        64'h02010913_08010993,
        64'h00050493_00010a93,
        64'hc61ff0ef_00010513,
        64'h00100613_e0010113,
        64'h04892583_d60ff0ef,
        64'h15050513_00001517,
        64'hdccff0ef_05412503,
        64'hd74ff0ef_34450513,
        64'h00001517_de0ff0ef,
        64'h05012503_d88ff0ef,
        64'h33850513_00001517,
        64'he54ff0ef_04813503,
        64'hd9cff0ef_32c50513,
        64'h00001517_e68ff0ef,
        64'h02013503_db0ff0ef,
        64'h33050513_00001517,
        64'he7cff0ef_01813503,
        64'hdc4ff0ef_32c50513,
        64'h00001517_e30ff0ef,
        64'h01412503_dd8ff0ef,
        64'h33050513_00001517,
        64'he44ff0ef_01012503,
        64'hdecff0ef_33450513,
        64'h00001517_e58ff0ef,
        64'h00c12503_e00ff0ef,
        64'h33850513_00001517,
        64'he6cff0ef_00812503,
        64'he14ff0ef_33c50513,
        64'h00001517_ee0ff0ef,
        64'h00013503_e28ff0ef,
        64'h34050513_00001517,
        64'he34ff0ef_32c50513,
        64'h00001517_f69ff06f,
        64'hffe00493_e48ff0ef,
        64'h23850513_00001517,
        64'hf14ff0ef_00048513,
        64'he5cff0ef_33c50513,
        64'h00001517_e68ff0ef,
        64'h33050513_00001517,
        64'h02050c63_00050493,
        64'h00010913_d95ff0ef,
        64'h00010513_00100593,
        64'h00100613_e0010113,
        64'he94ff0ef_34450513,
        64'h00001517_00008067,
        64'h06010113_00813c83,
        64'h01013c03_01813b83,
        64'h02013b03_02813a83,
        64'h03013a03_03813983,
        64'h04013903_04813483,
        64'h05013403_00048513,
        64'h05813083_fa040113,
        64'hfff00493_ee0ff0ef,
        64'h36850513_00001517,
        64'h04050863_d19ff0ef,
        64'h00050b13_06010413,
        64'h01913423_01813823,
        64'h01713c23_03513423,
        64'h03413823_03313c23,
        64'h05213023_04913423,
        64'h04113c23_03613023,
        64'h04813823_fa010113,
        64'hf85ff06f_ffe00413,
        64'h00008067_0d010113,
        64'h08813b83_09013b03,
        64'h09813a83_0a013a03,
        64'h0a813983_0b013903,
        64'h0b813483_0c013403,
        64'h0c813083_00040513,
        64'hfff00413_f68ff0ef,
        64'h3c850513_00001517,
        64'hb09ff0ef_b0dff0ef,
        64'hb11ff0ef_b15ff0ef,
        64'hb19ff0ef_b1dff0ef,
        64'hb21ff0ef_b25ff0ef,
        64'h0340006f_b2dff0ef,
        64'hb39ff0ef_00c00513,
        64'h00000593_00100613,
        64'h00000413_f73046e3,
        64'h20048493_fff98993,
        64'hfbcff0ef_43c50513,
        64'h00001517_00079863,
        64'h0369e7b3_0a891063,
        64'h03045413_0009091b,
        64'h03041413_00a46433,
        64'hb79ff0ef_03045413,
        64'h03051413_0085151b,
        64'hb89ff0ef_fc9412e3,
        64'h04040413_ff7a12e3,
        64'h00050913_ec1ff0ef,
        64'h0ff5f593_001a0a13,
        64'h00090513_0007c583,
        64'h014407b3_04000b93,
        64'h00000a13_b05ff0ef,
        64'h00010513_04000593,
        64'h00040613_00000913,
        64'hff551ee3_bd5ff0ef,
        64'he0048413_3e800b13,
        64'h0fe00a93_0c051063,
        64'h20048493_bf5ff0ef,
        64'h01200513_00040593,
        64'h0ff67613_00166613,
        64'h0015161b_f01ff0ef,
        64'h0ff47593_f09ff0ef,
        64'h0ff5f593_0084559b,
        64'hf15ff0ef_0ff5f593,
        64'h0104559b_f21ff0ef,
        64'h00000513_0184559b,
        64'hfee79ae3_00178793,
        64'h00c68023_00f106b3,
        64'h08000713_fff00613,
        64'h00000793_0209d993,
        64'h00058413_00050493,
        64'h09713423_09613823,
        64'h09513c23_0b413023,
        64'h0b213823_0c113423,
        64'h0a913c23_0c813023,
        64'h02061993_0b313423,
        64'hf3010113_00008067,
        64'h03055513_03051513,
        64'h00f54533_00e7f7b3,
        64'h0057979b_fe070713,
        64'h00002737_0107d79b,
        64'h0105179b_4105551b,
        64'h0105151b_00a5c533,
        64'h00c59513_00b545b3,
        64'h00f57513_0045d51b,
        64'h00b545b3_03055513,
        64'h03051513_00f56533,
        64'h00851513_0085579b,
        64'h00008067_07f57513,
        64'h00b54533_00451593,
        64'h00b54533_0ff57513,
        64'h00f54533_0045d51b,
        64'h0075d79b_00b575b3,
        64'h00008067_01010113,
        64'h00078513_00013403,
        64'h00813083_ffd00793,
        64'h00051463_00000793,
        64'hf5dff0ef_00050a63,
        64'hffe00793_e99ff0ef,
        64'h02050063_fff00793,
        64'he2dff0ef_fe041ce3,
        64'hd49ff0ef_fff4041b,
        64'h00a00413_9c1ff0ef,
        64'h60850513_00001517,
        64'hb2dff0ef_00813023,
        64'h00113423_ff010113,
        64'h00008067_02010113,
        64'h00153513_00813483,
        64'h01013403_01813083,
        64'h0004051b_fc940ae3,
        64'hd91ff0ef_e29ff0ef,
        64'h64050513_00001517,
        64'h00050593_00050413,
        64'hdb1ff0ef_02900513,
        64'h400005b7_07700613,
        64'hf9dff0ef_00100493,
        64'h00813823_00113c23,
        64'h00913423_fe010113,
        64'h00008067_01010113,
        64'h00153513_fff50513,
        64'h00013403_00813083,
        64'h0004051b_e81ff0ef,
        64'h69450513_00040593,
        64'h00001517_dfdff0ef,
        64'h00050413_e0dff0ef,
        64'h00813023_00113423,
        64'h03700513_00000593,
        64'h06500613_ff010113,
        64'h00008067_02010113,
        64'h00013903_00813483,
        64'h01013403_01813083,
        64'h00153513_f5650513,
        64'h0004051b_01249863,
        64'h00f4f493_00f91c63,
        64'h00000513_00100793,
        64'he59ff0ef_e5dff0ef,
        64'h00050413_e65ff0ef,
        64'h00050493_e6dff0ef,
        64'he71ff0ef_e75ff0ef,
        64'h00050913_e85ff0ef,
        64'h01213023_00913423,
        64'h00813823_00113c23,
        64'h00800513_1aa00593,
        64'h08700613_fe010113,
        64'hfe5ff06f_00000513,
        64'h00008067_02010113,
        64'h00013903_00813483,
        64'h01013403_01813083,
        64'h00100513_f59ff0ef,
        64'h00100593_76450513,
        64'h00001517_fe9910e3,
        64'h02040a63_eddff0ef,
        64'h00050913_fff4041b,
        64'hef1ff0ef_00000513,
        64'h00000593_09500613,
        64'h00100493_71040413,
        64'h01213023_00113c23,
        64'h00913423_00002437,
        64'h00813823_fe010113,
        64'hb85ff06f_02010113,
        64'h77850513_00001517,
        64'h01813083_01013403,
        64'hcbdff0ef_00058513,
        64'h00813583_ba9ff0ef,
        64'h7c850513_00001517,
        64'hbb5ff0ef_00040513,
        64'hbbdff0ef_00b13423,
        64'h00113c23_7d450513,
        64'h00001517_00050413,
        64'h00813823_fe010113,
        64'h00008067_03010113,
        64'h01813483_02013403,
        64'h02813083_fe0416e3,
        64'hfff40413_0007d663,
        64'h4187d79b_0185179b,
        64'hf99ff0ef_e31ff0ef,
        64'h00060513_06400413,
        64'h00813603_e41ff0ef,
        64'h0ff47513_e49ff0ef,
        64'h0ff57513_0084551b,
        64'he55ff0ef_0ff57513,
        64'h0104551b_e61ff0ef,
        64'h0184551b_e69ff0ef,
        64'h0404e513_fddff0ef,
        64'h00050493_00058413,
        64'h00913c23_02813023,
        64'h00c13423_02113423,
        64'hfd010113_e91ff06f,
        64'h0ff00513_00008067,
        64'hfff00513_fadff06f,
        64'h00d70023_00178793,
        64'h00f60733_06c82683,
        64'hfc0712e3_00177713,
        64'h06452703_f91ff06f,
        64'h06e6a423_00178793,
        64'h00074703_00f50733,
        64'h00008067_00000513,
        64'h06e7a023_00600713,
        64'h06e7a823_fff00713,
        64'h200007b7_02b6ea63,
        64'h0007869b_20000837,
        64'h20000537_fe079ce3,
        64'h0017f793_06472783,
        64'h20000737_06e7a023,
        64'h200007b7_10600713,
        64'hfe079ce3_fff7879b,
        64'h00000013_03200793,
        64'h04b76e63_0007871b,
        64'h00000793_200006b7,
        64'h06e7a823_ffe00713,
        64'h200007b7_0ab7e663,
        64'h10000793_00008067,
        64'h02010113_00813483,
        64'h06e7a023_00600713,
        64'h06e7a823_01013403,
        64'h01813083_0ff47513,
        64'hfff00713_200007b7,
        64'hd55ff0ef_94450513,
        64'h00002517_e21ff0ef,
        64'h02055513_02051513,
        64'h0004a503_d71ff0ef,
        64'h96850513_00002517,
        64'h02079663_0017f793,
        64'h0004041b_0647a783,
        64'h06c7a403_fe071ae3,
        64'h00177713_06478493,
        64'h0647a703_06e7a023,
        64'h10600713_200007b7,
        64'hfe079ce3_fff7879b,
        64'h00000013_06400793,
        64'h06a7a423_06e7a823,
        64'hffe00713_00913423,
        64'h00813823_00113c23,
        64'h200007b7_fe010113,
        64'hdddff06f_02010113,
        64'h9c050513_00002517,
        64'h00813483_01813083,
        64'h01013403_06f42023,
        64'h00600793_e01ff0ef,
        64'h9f050513_00002517,
        64'hecdff0ef_02055513,
        64'h02049513_0004849b,
        64'he1dff0ef_9ec50513,
        64'h00002517_06442483,
        64'h06f42023_16600793,
        64'he35ff0ef_a2450513,
        64'h00002517_f01ff0ef,
        64'h02055513_02049513,
        64'h0004849b_e51ff0ef,
        64'ha2050513_00002517,
        64'h06442483_06f42023,
        64'h10400793_20000437,
        64'hfe079ce3_fff7879b,
        64'h00000013_00a00793,
        64'h04e7a023_00a00713,
        64'h200007b7_e89ff0ef,
        64'h00913423_00813823,
        64'h00113c23_a5850513,
        64'hfe010113_00002517,
        64'h00008067_0005051b,
        64'h00052503_00008067,
        64'h00b52023_00008067,
        64'h02010113_01813083,
        64'he65ff0ef_00914503,
        64'he6dff0ef_00814503,
        64'hf09ff0ef_00113c23,
        64'h00810593_fe010113,
        64'h00008067_03010113,
        64'h01013903_01813483,
        64'h02013403_02813083,
        64'hfc941ee3_ea1ff0ef,
        64'h00914503_ea9ff0ef,
        64'hff84041b_00814503,
        64'hf49ff0ef_0ff57513,
        64'h00810593_00895533,
        64'hff800493_03800413,
        64'h00050913_02113423,
        64'h01213823_00913c23,
        64'h02813023_fd010113,
        64'h00008067_03010113,
        64'h01013903_01813483,
        64'h02013403_02813083,
        64'hfc941ee3_f01ff0ef,
        64'h00914503_f09ff0ef,
        64'hff84041b_00814503,
        64'hfa9ff0ef_0ff57513,
        64'h00810593_0089553b,
        64'hff800493_01800413,
        64'h00050913_02113423,
        64'h01213823_00913c23,
        64'h02813023_fd010113,
        64'h00008067_00f58023,
        64'h0007c783_00e580a3,
        64'h00a787b3_00455513,
        64'h00074703_00e78733,
        64'h00f57713_d4478793,
        64'h00001797_fe1ff06f,
        64'h00140413_f79ff0ef,
        64'h00008067_01010113,
        64'h00013403_00813083,
        64'h00051a63_00044503,
        64'h00050413_00113423,
        64'h00813023_ff010113,
        64'h00008067_00e78823,
        64'h02000713_00e78423,
        64'hfc700713_00e78623,
        64'h00300713_00a78223,
        64'h0ff57513_00e78023,
        64'h0085551b_0ff57713,
        64'h00e78623_f8000713,
        64'h00078223_100007b7,
        64'h02b5553b_0045959b,
        64'h00008067_00a70023,
        64'hfe078ce3_0207f793,
        64'h01474783_10000737,
        64'h00008067_02057513,
        64'h0147c503_100007b7,
        64'h00008067_0ff57513,
        64'h00054503_00008067,
        64'h00b50023_00008067,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00048067_01f49493,
        64'h0010049b_fa458593,
        64'h00001597_f1402573,
        64'h0924a4af_00190913,
        64'h04048493_01a49493,
        64'h0210049b_ff2496e3,
        64'hf14024f3_0004a903,
        64'h04048493_01a49493,
        64'h0210049b_59d000ef,
        64'h01a11113_0210011b,
        64'h01249863_f1402973,
        64'h00000493_0924a4af,
        64'h00000913_04048493,
        64'h01a49493_0210049b
    };

    logic [$clog2(RomSize)-1:0] addr_q;

    always_ff @(posedge clk_i) begin
        if (req_i) begin
            addr_q <= addr_i[$clog2(RomSize)-1+3:3];
        end
    end

    // this prevents spurious Xes from propagating into
    // the speculative fetch stage of the core
    assign rdata_o = (addr_q < RomSize) ? mem[addr_q] : '0;
endmodule
